* NGSPICE file created from Gilbert_mixer.ext - technology: gf180mcuD

.subckt Gilbert_mixer I_bias_p I_bias_n V_out_p V_out_n V_LO V_LO_b RF_POS RF_NEG
X0 I_bias_p RF_POS a_n572_n259# a_n1768_n2977# nfet_03v3 ad=1.22p pd=3.22u as=1.22p ps=3.22u w=2u l=0.28u M=5
X1 V_out_p V_LO I_bias_p a_n1768_n2977# nfet_03v3 ad=2.44p pd=5.22u as=2.44p ps=5.22u w=4u l=0.28u M=5
X2 a_n1768_n2977# a_n1768_n2977# a_n1768_n2977# a_n1768_n2977# nfet_03v3 ad=4.56p pd=10.28u as=91.2p ps=0.21472m w=4u l=0.28u M=8
X3 V_out_n V_LO_b I_bias_n a_n1768_n2977# nfet_03v3 ad=2.44p pd=5.22u as=2.44p ps=5.22u w=4u l=0.28u M=5
X4 I_bias_n RF_NEG a_n572_n2107# a_n1768_n2977# nfet_03v3 ad=1.22p pd=3.22u as=1.22p ps=3.22u w=2u l=0.28u M=5
X5 I_bias_n V_LO V_out_p a_n1768_n2977# nfet_03v3 ad=2.44p pd=5.22u as=2.44p ps=5.22u w=4u l=0.28u M=5
X6 a_n1768_n2977# a_n1768_n2977# a_n1768_n2977# a_n1768_n2977# nfet_03v3 ad=2.28p pd=6.28u as=0 ps=0 w=2u l=0.28u M=4
X7 I_bias_p V_LO_b V_out_n a_n1768_n2977# nfet_03v3 ad=2.44p pd=5.22u as=4.56p ps=10.28u w=4u l=0.28u M=5
.ends

