magic
tech gf180mcuD
magscale 1 10
timestamp 1757884110
<< pwell >>
rect -1176 -4755 1176 4755
<< mvpsubdiff >>
rect -1152 4718 1152 4731
rect -1152 4672 -1036 4718
rect 1036 4672 1152 4718
rect -1152 4659 1152 4672
rect -1152 4615 -1080 4659
rect -1152 2543 -1139 4615
rect -1093 2543 -1080 4615
rect 1080 4615 1152 4659
rect -1152 2499 -1080 2543
rect 1080 2543 1093 4615
rect 1139 2543 1152 4615
rect 1080 2499 1152 2543
rect -1152 2486 1152 2499
rect -1152 2440 -1036 2486
rect 1036 2440 1152 2486
rect -1152 2427 1152 2440
rect -1152 2332 1152 2345
rect -1152 2286 -1036 2332
rect 1036 2286 1152 2332
rect -1152 2273 1152 2286
rect -1152 2229 -1080 2273
rect -1152 157 -1139 2229
rect -1093 157 -1080 2229
rect 1080 2229 1152 2273
rect -1152 113 -1080 157
rect 1080 157 1093 2229
rect 1139 157 1152 2229
rect 1080 113 1152 157
rect -1152 100 1152 113
rect -1152 54 -1036 100
rect 1036 54 1152 100
rect -1152 41 1152 54
rect -1152 -54 1152 -41
rect -1152 -100 -1036 -54
rect 1036 -100 1152 -54
rect -1152 -113 1152 -100
rect -1152 -157 -1080 -113
rect -1152 -2229 -1139 -157
rect -1093 -2229 -1080 -157
rect 1080 -157 1152 -113
rect -1152 -2273 -1080 -2229
rect 1080 -2229 1093 -157
rect 1139 -2229 1152 -157
rect 1080 -2273 1152 -2229
rect -1152 -2286 1152 -2273
rect -1152 -2332 -1036 -2286
rect 1036 -2332 1152 -2286
rect -1152 -2345 1152 -2332
rect -1152 -2440 1152 -2427
rect -1152 -2486 -1036 -2440
rect 1036 -2486 1152 -2440
rect -1152 -2499 1152 -2486
rect -1152 -2543 -1080 -2499
rect -1152 -4615 -1139 -2543
rect -1093 -4615 -1080 -2543
rect 1080 -2543 1152 -2499
rect -1152 -4659 -1080 -4615
rect 1080 -4615 1093 -2543
rect 1139 -4615 1152 -2543
rect 1080 -4659 1152 -4615
rect -1152 -4672 1152 -4659
rect -1152 -4718 -1036 -4672
rect 1036 -4718 1152 -4672
rect -1152 -4731 1152 -4718
<< mvpsubdiffcont >>
rect -1036 4672 1036 4718
rect -1139 2543 -1093 4615
rect 1093 2543 1139 4615
rect -1036 2440 1036 2486
rect -1036 2286 1036 2332
rect -1139 157 -1093 2229
rect 1093 157 1139 2229
rect -1036 54 1036 100
rect -1036 -100 1036 -54
rect -1139 -2229 -1093 -157
rect 1093 -2229 1139 -157
rect -1036 -2332 1036 -2286
rect -1036 -2486 1036 -2440
rect -1139 -4615 -1093 -2543
rect 1093 -4615 1139 -2543
rect -1036 -4718 1036 -4672
<< mvndiode >>
rect -1000 4566 1000 4579
rect -1000 2592 -987 4566
rect 987 2592 1000 4566
rect -1000 2579 1000 2592
rect -1000 2180 1000 2193
rect -1000 206 -987 2180
rect 987 206 1000 2180
rect -1000 193 1000 206
rect -1000 -206 1000 -193
rect -1000 -2180 -987 -206
rect 987 -2180 1000 -206
rect -1000 -2193 1000 -2180
rect -1000 -2592 1000 -2579
rect -1000 -4566 -987 -2592
rect 987 -4566 1000 -2592
rect -1000 -4579 1000 -4566
<< mvndiodec >>
rect -987 2592 987 4566
rect -987 206 987 2180
rect -987 -2180 987 -206
rect -987 -4566 987 -2592
<< metal1 >>
rect -1139 4672 -1036 4718
rect 1036 4672 1139 4718
rect -1139 4615 -1093 4672
rect 1093 4615 1139 4672
rect -998 2592 -987 4566
rect 987 2592 998 4566
rect -1139 2486 -1093 2543
rect 1093 2486 1139 2543
rect -1139 2440 -1036 2486
rect 1036 2440 1139 2486
rect -1139 2286 -1036 2332
rect 1036 2286 1139 2332
rect -1139 2229 -1093 2286
rect 1093 2229 1139 2286
rect -998 206 -987 2180
rect 987 206 998 2180
rect -1139 100 -1093 157
rect 1093 100 1139 157
rect -1139 54 -1036 100
rect 1036 54 1139 100
rect -1139 -100 -1036 -54
rect 1036 -100 1139 -54
rect -1139 -157 -1093 -100
rect 1093 -157 1139 -100
rect -998 -2180 -987 -206
rect 987 -2180 998 -206
rect -1139 -2286 -1093 -2229
rect 1093 -2286 1139 -2229
rect -1139 -2332 -1036 -2286
rect 1036 -2332 1139 -2286
rect -1139 -2486 -1036 -2440
rect 1036 -2486 1139 -2440
rect -1139 -2543 -1093 -2486
rect 1093 -2543 1139 -2486
rect -998 -4566 -987 -2592
rect 987 -4566 998 -2592
rect -1139 -4672 -1093 -4615
rect 1093 -4672 1139 -4615
rect -1139 -4718 -1036 -4672
rect 1036 -4718 1139 -4672
<< properties >>
string diode_nd2ps_06v0_9F7TZ3 parameters
string FIXED_BBOX -1116 2463 1116 4695
string gencell diode_nd2ps_06v0
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 1 ny 4 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 doverlap 0 full_metal 1 compatible {diode_nd2ps_03v3 diode_nd2ps_06v0}
<< end >>
