magic
tech gf180mcuD
magscale 1 10
timestamp 1755084777
<< error_p >>
rect -354 2033 -343 2079
rect -297 2033 -286 2044
rect -194 2033 -183 2079
rect -137 2033 -126 2044
rect -34 2033 -23 2079
rect 23 2033 34 2044
rect 126 2033 137 2079
rect 183 2033 194 2044
rect 286 2033 297 2079
rect 343 2033 354 2044
rect -400 -1998 -377 -1987
rect -263 -1998 -217 -1987
rect -103 -1998 -57 -1987
rect 57 -1998 103 -1987
rect 217 -1998 263 -1987
rect 377 -1998 400 -1987
rect -354 -2079 -343 -2033
rect -194 -2079 -183 -2033
rect -34 -2079 -23 -2033
rect 126 -2079 137 -2033
rect 286 -2079 297 -2033
<< pwell >>
rect -598 -2210 598 2210
<< nmos >>
rect -348 -2000 -292 2000
rect -188 -2000 -132 2000
rect -28 -2000 28 2000
rect 132 -2000 188 2000
rect 292 -2000 348 2000
<< ndiff >>
rect -436 1987 -348 2000
rect -436 -1987 -423 1987
rect -377 -1987 -348 1987
rect -436 -2000 -348 -1987
rect -292 1987 -188 2000
rect -292 -1987 -263 1987
rect -217 -1987 -188 1987
rect -292 -2000 -188 -1987
rect -132 1987 -28 2000
rect -132 -1987 -103 1987
rect -57 -1987 -28 1987
rect -132 -2000 -28 -1987
rect 28 1987 132 2000
rect 28 -1987 57 1987
rect 103 -1987 132 1987
rect 28 -2000 132 -1987
rect 188 1987 292 2000
rect 188 -1987 217 1987
rect 263 -1987 292 1987
rect 188 -2000 292 -1987
rect 348 1987 436 2000
rect 348 -1987 377 1987
rect 423 -1987 436 1987
rect 348 -2000 436 -1987
<< ndiffc >>
rect -423 -1987 -377 1987
rect -263 -1987 -217 1987
rect -103 -1987 -57 1987
rect 57 -1987 103 1987
rect 217 -1987 263 1987
rect 377 -1987 423 1987
<< psubdiff >>
rect -574 2114 574 2186
rect -574 2070 -502 2114
rect -574 -2070 -561 2070
rect -515 -2070 -502 2070
rect 502 2070 574 2114
rect -574 -2114 -502 -2070
rect 502 -2070 515 2070
rect 561 -2070 574 2070
rect 502 -2114 574 -2070
rect -574 -2186 574 -2114
<< psubdiffcont >>
rect -561 -2070 -515 2070
rect 515 -2070 561 2070
<< polysilicon >>
rect -356 2079 -284 2092
rect -356 2033 -343 2079
rect -297 2033 -284 2079
rect -356 2020 -284 2033
rect -196 2079 -124 2092
rect -196 2033 -183 2079
rect -137 2033 -124 2079
rect -196 2020 -124 2033
rect -36 2079 36 2092
rect -36 2033 -23 2079
rect 23 2033 36 2079
rect -36 2020 36 2033
rect 124 2079 196 2092
rect 124 2033 137 2079
rect 183 2033 196 2079
rect 124 2020 196 2033
rect 284 2079 356 2092
rect 284 2033 297 2079
rect 343 2033 356 2079
rect 284 2020 356 2033
rect -348 2000 -292 2020
rect -188 2000 -132 2020
rect -28 2000 28 2020
rect 132 2000 188 2020
rect 292 2000 348 2020
rect -348 -2020 -292 -2000
rect -188 -2020 -132 -2000
rect -28 -2020 28 -2000
rect 132 -2020 188 -2000
rect 292 -2020 348 -2000
rect -356 -2033 -284 -2020
rect -356 -2079 -343 -2033
rect -297 -2079 -284 -2033
rect -356 -2092 -284 -2079
rect -196 -2033 -124 -2020
rect -196 -2079 -183 -2033
rect -137 -2079 -124 -2033
rect -196 -2092 -124 -2079
rect -36 -2033 36 -2020
rect -36 -2079 -23 -2033
rect 23 -2079 36 -2033
rect -36 -2092 36 -2079
rect 124 -2033 196 -2020
rect 124 -2079 137 -2033
rect 183 -2079 196 -2033
rect 124 -2092 196 -2079
rect 284 -2033 356 -2020
rect 284 -2079 297 -2033
rect 343 -2079 356 -2033
rect 284 -2092 356 -2079
<< polycontact >>
rect -343 2033 -297 2079
rect -183 2033 -137 2079
rect -23 2033 23 2079
rect 137 2033 183 2079
rect 297 2033 343 2079
rect -343 -2079 -297 -2033
rect -183 -2079 -137 -2033
rect -23 -2079 23 -2033
rect 137 -2079 183 -2033
rect 297 -2079 343 -2033
<< metal1 >>
rect -561 2127 561 2173
rect -561 2070 -515 2127
rect -354 2033 -343 2079
rect -297 2033 -286 2079
rect -194 2033 -183 2079
rect -137 2033 -126 2079
rect -34 2033 -23 2079
rect 23 2033 34 2079
rect 126 2033 137 2079
rect 183 2033 194 2079
rect 286 2033 297 2079
rect 343 2033 354 2079
rect 515 2070 561 2127
rect -423 1987 -377 1998
rect -423 -1998 -377 -1987
rect -263 1987 -217 1998
rect -263 -1998 -217 -1987
rect -103 1987 -57 1998
rect -103 -1998 -57 -1987
rect 57 1987 103 1998
rect 57 -1998 103 -1987
rect 217 1987 263 1998
rect 217 -1998 263 -1987
rect 377 1987 423 1998
rect 377 -1998 423 -1987
rect -561 -2127 -515 -2070
rect -354 -2079 -343 -2033
rect -297 -2079 -286 -2033
rect -194 -2079 -183 -2033
rect -137 -2079 -126 -2033
rect -34 -2079 -23 -2033
rect 23 -2079 34 -2033
rect 126 -2079 137 -2033
rect 183 -2079 194 -2033
rect 286 -2079 297 -2033
rect 343 -2079 354 -2033
rect 515 -2127 561 -2070
rect -561 -2173 561 -2127
<< properties >>
string FIXED_BBOX -538 -2150 538 2150
string gencell nfet_03v3
string library gf180mcu
string parameters w 20.0 l 0.28 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
