** sch_path: /foss/designs/Chipathon_2025_gLayout/src/design_tb/Gilbert_cell_tb_IIP3.sch
**.subckt Gilbert_cell_tb_IIP3 V_LO V_LO_b V_RF V_RF_b V_out_p V_out_n
*.ipin V_LO
*.ipin V_LO_b
*.ipin V_RF
*.ipin V_RF_b
*.opin V_out_p
*.opin V_out_n
V_PWR VDD GND 3.3
.save i(v_pwr)
V_LO V_LO GND pulse(0 1.5 0 1p 1p 0.25n 0.5n)
.save i(v_lo)
V_LO_b V_LO_b GND pulse(0 1.5 0 1p 1p 0.25n 0.5n)
.save i(v_lo_b)
V_RF_tone_1 net2 GND sin( 1 1 1 0 )
.save i(v_rf_tone_1)
V_RF_b_tone_1 net1 GND sin( 1 1 1 0 0 180 )
.save i(v_rf_b_tone_1)
xGilbert_mixer VDD V_out_n V_out_p V_LO V_LO_b V_RF_b V_RF I_bias_pos I_bias_neg GND Gilbert_cell_no_hierarchy
I0 I_bias_pos GND 50u
I1 I_bias_neg GND 50u
V_RF_tone_2 V_RF net2 sin( 1 1 1 0 )
.save i(v_rf_tone_2)
V_RF_b_tone_2 V_RF_b net1 sin( 1 1 1 0 0 180 )
.save i(v_rf_b_tone_2)
**** begin user architecture code

.include /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /usr/local/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical




* let sets vectors to a plot, while set sets a variable, globally accessible in .control
.control

    * Set frequency and amplitude variables to proper values from within the control sequence
    set freq_lo = 100Meg
    set cm_lo = 1.6
    set amp_lo = 0.4

    set cm_rf  = 0.6
    set freq_rf_tone_1 = 89.3Meg
    set freq_rf_tone_2 = 89.4Meg
    set amp_rf  = 0.1

    * set the parameters to the voltage sources
    alter @V_LO[sin] = [ $cm_lo $amp_lo $freq_lo 0 ]
    alter @V_LO_b[sin] = [ $cm_lo $amp_lo $freq_lo 0 0 180 ]
    alter @V_RF_tone_1[sin] = [ $cm_rf $amp_rf $freq_rf_tone_1 0 ]
    alter @V_RF_b_tone_1[sin] = [ $cm_rf $amp_rf $freq_rf_tone_1 0 0 180 ]
    alter @V_RF_tone_2[sin] = [ $cm_rf $amp_rf $freq_rf_tone_2 0 ]
    alter @V_RF_b_tone_2[sin] = [ $cm_rf $amp_rf $freq_rf_tone_2 0 0 180 ]

    save all

    * operating point
    * op
    * show


    * Transient analysis to observe mixing operation
    tran 0.1p 10u
    write Gilbert_cell_tb_IIP3_sim.raw

    set appendwrite

    * Calculate differential output for conversion gain measurement
    let v_out_diff = v(v_out_p)-v(v_out_n)
    let v_rf_diff = v(v_rf)-v(v_rf_b)
    let v_lo_diff = v(v_lo)-v(v_lo_b)


    * Extract IF component at 100MHz using FFT
    linearize v_out_diff v_rf_diff v_lo_diff
    let time_step = 1e-12
    let sample_freq = 1/time_step
    let npts = length(v_out_diff)
    let freq_res = sample_freq/npts

    fft v_out_diff v_rf_diff v_lo_diff
    * Find frequency bins

    * print everything, sanity check
    * set     ; print all available global (?) variables (?)
    * setplot ; print all plots
    * display ; print variables available in current plot

    let freq_res = tran2.freq_res
    let freq_if_1 = abs( $freq_lo - $freq_rf_tone_1)
    let freq_if_2 = abs( $freq_lo - $freq_rf_tone_2)

    let if_bin_1 = floor( freq_if_1/freq_res )
    let if_bin_2 = floor( freq_if_2/freq_res )
    let rf_bin_1 = floor( $freq_rf_tone_1/freq_res )
    let rf_bin_2 = floor( $freq_rf_tone_2/freq_res )

    * Measure conversion gain (power gain from RF to IF)
    * let rf_tone_1_mag = abs(v_rf_tone_1_diff[rf_bin_1])
    * let rf_tone_2_mag = abs(v_rf_tone_2_diff[rf_bin_2])
    * let if_mag = abs(v_out_diff[if_bin])
    * let conversion_gain_db = 20*log10(if_mag/rf_mag)
    * print conversion_gain_db

    write Gilbert_cell_tb_IIP3_sim.raw

.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/Chipathon_2025_gLayout/src/design_xsch/Gilbert_cell_no_hierarchy.sym # of pins=10
** sym_path: /foss/designs/Chipathon_2025_gLayout/src/design_xsch/Gilbert_cell_no_hierarchy.sym
** sch_path: /foss/designs/Chipathon_2025_gLayout/src/design_xsch/Gilbert_cell_no_hierarchy.sch
.subckt Gilbert_cell_no_hierarchy VDD V_out_p V_out_n V_LO V_LO_b V_RF V_RF_b I_bias_pos I_bias_neg VSS
*.ipin V_LO
*.ipin V_LO_b
*.ipin V_RF
*.ipin V_RF_b
*.opin V_out_p
*.opin V_out_n
*.iopin I_bias_neg
*.iopin I_bias_pos
*.iopin VDD
*.iopin VSS
R1 VDD V_out_p 6K m=1
R2 VDD V_out_n 6K m=1
XM_dp_lo_pos V_out_p V_LO rf_diff_pair_pos_input VSS nfet_03v3 L=0.28u W=20u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM_dp_lo_neg V_out_n V_LO_b rf_diff_pair_pos_input VSS nfet_03v3 L=0.28u W=20u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM_dp_lo_b_pos V_out_p V_LO_b rf_diff_pair_neg_input VSS nfet_03v3 L=0.28u W=20u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM_dp_lo_b_neg V_out_n V_LO rf_diff_pair_neg_input VSS nfet_03v3 L=0.28u W=20u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM_rf_pos rf_diff_pair_pos_input V_RF I_bias_pos VSS nfet_03v3 L=0.28u W=10u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM_rf_neg rf_diff_pair_neg_input V_RF_b I_bias_neg VSS nfet_03v3 L=0.28u W=10u nf=5 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
R7 I_bias_pos I_bias_neg 2K m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
