magic
tech gf180mcuD
magscale 1 10
timestamp 1757933240
<< metal1 >>
rect -7502 6590 2533 7015
rect -7502 6264 -6544 6590
rect 2161 6264 2533 6590
rect -7502 6210 2533 6264
rect 2218 5926 2302 5928
rect -6653 5836 -6638 5926
rect 2279 5836 2302 5926
rect 2218 5830 2302 5836
rect -6289 3802 -6279 4386
rect -4938 3802 -4928 4386
rect -4069 3823 -4059 4407
rect -2718 3823 -2708 4407
rect -1849 3809 -1839 4393
rect -498 3809 -488 4393
rect 378 3823 388 4407
rect 1729 3823 1739 4407
rect -7110 2210 2650 2400
rect -7110 30 -6660 2210
rect -6282 1397 -6272 1981
rect -4931 1397 -4921 1981
rect -4065 1397 -4055 1981
rect -2714 1397 -2704 1981
rect -1848 1418 -1838 2002
rect -497 1418 -487 2002
rect 369 1408 379 1992
rect 1720 1408 1730 1992
rect 2200 30 2650 2210
rect -7110 -990 2650 30
<< via1 >>
rect -6544 6264 2161 6590
rect -6638 5836 2279 5926
rect -6279 3802 -4938 4386
rect -4059 3823 -2718 4407
rect -1839 3809 -498 4393
rect 388 3823 1729 4407
rect -6272 1397 -4931 1981
rect -4055 1397 -2714 1981
rect -1838 1418 -497 2002
rect 379 1408 1720 1992
<< metal2 >>
rect -6662 6590 2310 6721
rect -6662 6264 -6544 6590
rect 2161 6264 2310 6590
rect -6662 6158 2310 6264
rect -6660 5926 2309 6158
rect -6660 5836 -6638 5926
rect 2279 5836 2309 5926
rect -6660 5823 2309 5836
rect -6304 4386 -4898 4441
rect -6304 3802 -6279 4386
rect -4938 3802 -4898 4386
rect -6304 3175 -4898 3802
rect -4084 4407 -2678 4450
rect -4084 3823 -4059 4407
rect -2718 3823 -2678 4407
rect -4084 3175 -2678 3823
rect -1865 4393 -459 4448
rect -1865 3809 -1839 4393
rect -498 3809 -459 4393
rect -1865 3175 -459 3809
rect 350 4407 1756 4462
rect 350 3823 388 4407
rect 1729 3823 1756 4407
rect 350 3175 1756 3823
rect -7396 2610 3274 3175
rect -6304 1981 -4898 2610
rect -4084 2510 -2677 2610
rect -6304 1397 -6272 1981
rect -4931 1397 -4898 1981
rect -6304 1360 -4898 1397
rect -4083 1981 -2677 2510
rect -4083 1397 -4055 1981
rect -2714 1397 -2677 1981
rect -4083 1365 -2677 1397
rect -1865 2002 -459 2610
rect 350 2522 1757 2610
rect -1865 1418 -1838 2002
rect -497 1418 -459 2002
rect -1865 1382 -459 1418
rect 351 1992 1757 2522
rect 351 1408 379 1992
rect 1720 1408 1757 1992
rect 351 1375 1757 1408
use diode_nd2ps_06v0_MV3SZ3  diode_nd2ps_06v0_MV3SZ3_0
timestamp 1757928106
transform 1 0 -2232 0 1 1116
box -4524 -1176 4524 1176
use diode_pd2nw_06v0_5DG9HC  diode_pd2nw_06v0_5DG9HC_0
timestamp 1757928106
transform 1 0 -2174 0 1 4732
box -4676 -1352 4676 1352
use ppolyf_u_4VJXJK  ppolyf_u_4VJXJK_0
timestamp 1757928106
transform 0 1 4548 -1 0 3036
box -1816 -718 1816 718
<< labels >>
rlabel metal1 -7010 -610 -7010 -610 1 VSS
port 0 n
rlabel metal2 -7307 2849 -7307 2849 1 to_gate
port 1 n
rlabel metal1 -7397 6678 -7397 6678 1 VDD
port 2 n
<< end >>
