magic
tech gf180mcuD
magscale 1 10
timestamp 1758010554
<< metal1 >>
rect -6440 12150 7520 12240
rect -6440 12140 5110 12150
rect -6440 11530 -6410 12140
rect 2510 11530 5110 12140
rect -6440 11450 5110 11530
rect 4140 11448 5110 11450
rect -8460 9820 -6510 9850
rect -8460 -4800 -8390 9820
rect -6880 7290 -6510 9820
rect -6420 9710 -6370 9720
rect 2490 9710 2540 9720
rect -6420 9620 -6410 9710
rect 2507 9620 2540 9710
rect -6420 9610 -6370 9620
rect 2490 9610 2540 9620
rect -5940 8480 -4580 8490
rect -5940 8316 -5930 8480
rect -5943 7732 -5930 8316
rect -5940 7730 -5930 7732
rect -4590 7730 -4580 8480
rect 680 8470 2040 8480
rect -3720 8460 -2360 8470
rect -3720 8297 -3710 8460
rect -5940 7720 -4580 7730
rect -3726 7713 -3710 8297
rect -3720 7710 -3710 7713
rect -2370 7710 -2360 8460
rect -1500 8460 -140 8470
rect -1500 8293 -1490 8460
rect -3720 7700 -2360 7710
rect -1501 7710 -1490 8293
rect -150 7710 -140 8460
rect 680 7720 690 8470
rect 2030 8307 2040 8470
rect 2030 7723 2041 8307
rect 2030 7720 2040 7723
rect 680 7710 2040 7720
rect -1501 7709 -140 7710
rect -1500 7700 -140 7709
rect 2620 7290 2950 9850
rect 4160 7410 5110 11448
rect -6880 -1620 2950 7290
rect -6880 -1650 -6360 -1620
rect 2500 -1650 2950 -1620
rect 4170 7090 5110 7410
rect 6620 7090 7520 12150
rect 4170 6880 7520 7090
rect 4170 -1340 4630 6880
rect 4680 6760 4810 6770
rect 4680 -1230 4690 6760
rect 4800 -1230 4810 6760
rect 4680 -1240 4810 -1230
rect 6880 6760 7010 6770
rect 6880 -1230 6890 6760
rect 7000 -1230 7010 6760
rect 6880 -1240 7010 -1230
rect 7070 -1340 7520 6880
rect -6880 -3810 -6358 -1650
rect -5940 -1829 -4580 -1820
rect -3720 -1829 -2360 -1820
rect -5942 -1830 -4580 -1829
rect -5942 -2413 -5930 -1830
rect -5940 -2580 -5930 -2413
rect -4590 -2580 -4580 -1830
rect -3725 -1830 -2360 -1829
rect -3725 -2413 -3710 -1830
rect -5940 -2590 -4580 -2580
rect -3720 -2580 -3710 -2413
rect -2370 -2580 -2360 -1830
rect -3720 -2590 -2360 -2580
rect -1500 -1826 -140 -1820
rect 680 -1826 2040 -1820
rect -1500 -1830 -139 -1826
rect -1500 -2580 -1490 -1830
rect -150 -2410 -139 -1830
rect 680 -1830 2041 -1826
rect -150 -2580 -140 -2410
rect -1500 -2590 -140 -2580
rect 680 -2580 690 -1830
rect 2030 -2410 2041 -1830
rect 2500 -1880 2952 -1650
rect 2030 -2580 2040 -2410
rect 680 -2590 2040 -2580
rect 2502 -3810 2952 -1880
rect 4170 -2070 7520 -1340
rect -6880 -4800 2952 -3810
rect -8460 -4830 2952 -4800
<< via1 >>
rect -6410 11530 2510 12140
rect -8390 -4800 -6880 9820
rect -6410 9620 2507 9710
rect -5930 7730 -4590 8480
rect -3710 7710 -2370 8460
rect -1490 7710 -150 8460
rect 690 7720 2030 8470
rect 5110 7090 6620 12150
rect 4690 -1230 4800 6760
rect 6890 -1230 7000 6760
rect -5930 -2580 -4590 -1830
rect -3710 -2580 -2370 -1830
rect -1490 -2580 -150 -1830
rect 690 -2580 2030 -1830
<< metal2 >>
rect -6440 12140 2540 12190
rect -6440 11530 -6410 12140
rect 2510 11530 2540 12140
rect -6440 11520 2540 11530
rect -6433 11388 2540 11520
rect -6431 11120 2540 11388
rect -8400 9820 -6870 9830
rect -8400 -4800 -8390 9820
rect -6880 -4800 -6870 9820
rect -6430 9710 2540 11120
rect -6430 9620 -6410 9710
rect 2507 9620 2540 9710
rect -6430 9600 2540 9620
rect 5100 12150 6630 12160
rect -5940 8490 -4580 8500
rect 680 8480 2040 8490
rect -5950 7732 -5940 8330
rect -3720 8470 -2360 8480
rect -4580 7732 -4570 8330
rect -3730 7713 -3720 8330
rect -5940 7700 -4580 7710
rect -1500 8470 -140 8480
rect -2360 7713 -2350 8330
rect -1510 7709 -1500 8330
rect -3720 7680 -2360 7690
rect -140 7709 -130 8330
rect 670 7723 680 8320
rect 2040 7723 2050 8320
rect 680 7690 2040 7700
rect -1500 7680 -140 7690
rect 5100 7090 5110 12150
rect 6620 7090 6630 12150
rect 5100 7080 6630 7090
rect 4620 6760 4810 6770
rect 4620 -1230 4640 6760
rect 4800 -1230 4810 6760
rect 4620 -1240 4810 -1230
rect 6880 6760 7050 6770
rect 6880 -1230 6890 6760
rect 6880 -1240 7050 -1230
rect -5940 -1810 -4580 -1800
rect -5950 -2420 -5940 -1829
rect -3720 -1810 -2360 -1800
rect -4580 -2420 -4570 -1829
rect -3730 -2420 -3720 -1829
rect -1500 -1810 -140 -1800
rect -5940 -2600 -4580 -2590
rect -2360 -2420 -2350 -1829
rect -1510 -2420 -1500 -1826
rect 680 -1810 2040 -1800
rect -3720 -2600 -2360 -2590
rect -140 -2420 -130 -1826
rect 670 -2430 680 -1826
rect -1500 -2600 -140 -2590
rect 2040 -2430 2050 -1826
rect 680 -2600 2040 -2590
rect -8400 -4810 -6870 -4800
<< via2 >>
rect -5940 8480 -4580 8490
rect -5940 7730 -5930 8480
rect -5930 7730 -4590 8480
rect -4590 7730 -4580 8480
rect -3720 8460 -2360 8470
rect -5940 7710 -4580 7730
rect -3720 7710 -3710 8460
rect -3710 7710 -2370 8460
rect -2370 7710 -2360 8460
rect -1500 8460 -140 8470
rect -3720 7690 -2360 7710
rect -1500 7710 -1490 8460
rect -1490 7710 -150 8460
rect -150 7710 -140 8460
rect 680 8470 2040 8480
rect -1500 7690 -140 7710
rect 680 7720 690 8470
rect 690 7720 2030 8470
rect 2030 7720 2040 8470
rect 680 7700 2040 7720
rect 4640 -1230 4690 6760
rect 4690 -1230 4800 6760
rect 6890 -1230 7000 6760
rect 7000 -1230 7050 6760
rect -5940 -1830 -4580 -1810
rect -5940 -2580 -5930 -1830
rect -5930 -2580 -4590 -1830
rect -4590 -2580 -4580 -1830
rect -3720 -1830 -2360 -1810
rect -5940 -2590 -4580 -2580
rect -3720 -2580 -3710 -1830
rect -3710 -2580 -2370 -1830
rect -2370 -2580 -2360 -1830
rect -1500 -1830 -140 -1810
rect -3720 -2590 -2360 -2580
rect -1500 -2580 -1490 -1830
rect -1490 -2580 -150 -1830
rect -150 -2580 -140 -1830
rect 680 -1830 2040 -1810
rect -1500 -2590 -140 -2580
rect 680 -2580 690 -1830
rect 690 -2580 2030 -1830
rect 2030 -2580 2040 -1830
rect 680 -2590 2040 -2580
<< metal3 >>
rect -5950 7710 -5940 8490
rect -4580 7710 -4570 8490
rect -5950 6760 -4570 7710
rect -3730 7690 -3720 8470
rect -2360 7690 -2350 8470
rect -3730 6760 -2350 7690
rect -1510 7690 -1500 8470
rect -140 7690 -130 8470
rect -1510 6760 -130 7690
rect 670 7700 680 8480
rect 2040 7700 2050 8480
rect 670 6760 2050 7700
rect 6880 6760 7760 6770
rect -8460 -1230 4640 6760
rect 4800 -1230 4810 6760
rect 6880 -1230 6890 6760
rect 7050 -1230 7760 6760
rect -8460 -1240 4690 -1230
rect 6880 -1240 7760 -1230
rect -5950 -1810 -4570 -1240
rect -5950 -2590 -5940 -1810
rect -4580 -2590 -4570 -1810
rect -3730 -1810 -2350 -1240
rect -3730 -2590 -3720 -1810
rect -2360 -2590 -2350 -1810
rect -1510 -1810 -130 -1240
rect -1510 -2590 -1500 -1810
rect -140 -2590 -130 -1810
rect 670 -1810 2050 -1240
rect 670 -2590 680 -1810
rect 2040 -2590 2050 -1810
use diode_nd2ps_06v0_MV3SZ3  diode_nd2ps_06v0_MV3SZ3_0
timestamp 1757961865
transform 1 0 -1916 0 1 -2714
box -4524 -1176 4524 1176
use diode_pd2nw_06v0_5DG9HC  diode_pd2nw_06v0_5DG9HC_0
timestamp 1757961865
transform 1 0 -1944 0 1 8542
box -4676 -1352 4676 1352
use ppolyf_u_9H3LNU  ppolyf_u_9H3LNU_0
timestamp 1757961865
transform 0 1 5848 -1 0 2766
box -4216 -1318 4216 1318
<< labels >>
rlabel metal1 -6708 -4450 -6708 -4450 1 VSS
port 3 n
rlabel metal3 -7870 3090 -7870 3090 1 to_gate
port 1 n
rlabel metal3 7600 2930 7600 2930 1 ASIG5V
port 0 n
rlabel via1 5760 11670 5760 11670 1 VDD
port 2 n
<< end >>
