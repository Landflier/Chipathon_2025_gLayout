* NGSPICE file created from pmos_Cmirror_with_decap_layout.ext - technology: gf180mcuD

.subckt Unnamed_ad0e3c17 m4_n620_n620# m4_n500_n500#
X0 m4_n500_n500# m4_n620_n620# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt cmirror_interdigitized a_n1022_n50# w_n2172_n840# a_n1856_n470#
X0 w_n2172_n840# a_n1856_n470# a_n1022_n50# w_n2172_n840# pfet_03v3 ad=0.305p pd=1.72u as=0.305p ps=1.72u w=0.5u l=0.28u M=8
X1 w_n2172_n840# a_n1856_n470# a_n1856_n470# w_n2172_n840# pfet_03v3 ad=0.305p pd=1.72u as=0.305p ps=1.72u w=0.5u l=0.28u M=4
.ends

.subckt pmos_Cmirror_with_decap_layout I_BIAS I_OUT VDD
XUnnamed_ad0e3c17_0 I_BIAS VDD Unnamed_ad0e3c17
Xcmirror_interdigitized_0 I_OUT VDD I_BIAS cmirror_interdigitized
.ends

