magic
tech gf180mcuD
magscale 1 10
timestamp 1757928606
<< metal1 >>
rect -7110 2210 2650 2400
rect -7110 30 -6660 2210
rect -6282 1397 -6272 1981
rect -4931 1397 -4921 1981
rect -4065 1397 -4055 1981
rect -2714 1397 -2704 1981
rect -1848 1418 -1838 2002
rect -497 1418 -487 2002
rect 369 1408 379 1992
rect 1720 1408 1730 1992
rect 2200 30 2650 2210
rect -7110 -990 2650 30
<< via1 >>
rect -6272 1397 -4931 1981
rect -4055 1397 -2714 1981
rect -1838 1418 -497 2002
rect 379 1408 1720 1992
<< metal2 >>
rect -7396 2610 3274 3175
rect -6304 1981 -4898 2610
rect -6304 1397 -6272 1981
rect -4931 1397 -4898 1981
rect -6304 1360 -4898 1397
rect -4083 1981 -2677 2610
rect -4083 1397 -4055 1981
rect -2714 1397 -2677 1981
rect -4083 1365 -2677 1397
rect -1865 2002 -459 2610
rect -1865 1418 -1838 2002
rect -497 1418 -459 2002
rect -1865 1382 -459 1418
rect 351 1992 1757 2610
rect 351 1408 379 1992
rect 1720 1408 1757 1992
rect 351 1375 1757 1408
use diode_nd2ps_06v0_MV3SZ3  diode_nd2ps_06v0_MV3SZ3_0
timestamp 1757928106
transform 1 0 -2232 0 1 1116
box -4524 -1176 4524 1176
use diode_pd2nw_06v0_5DG9HC  diode_pd2nw_06v0_5DG9HC_0
timestamp 1757928106
transform 1 0 -2174 0 1 4732
box -4676 -1352 4676 1352
use ppolyf_u_4VJXJK  ppolyf_u_4VJXJK_0
timestamp 1757928106
transform 0 1 4548 -1 0 3036
box -1816 -718 1816 718
<< labels >>
rlabel metal1 -7010 -610 -7010 -610 1 VSS
port 0 n
rlabel metal2 -7307 2849 -7307 2849 1 to_gate
port 1 n
<< end >>
