** sch_path: /home/vasil/Downloads/SSCS_PICO_2025/src/python/Gilbert_mixer_intedigited/Gilbert_cell_hierarchal_mixing_stage.sch
.subckt Gilbert_cell_hierarchal_mixing_stage V_out_n V_out_p V_LO V_LO_b V_RF V_RF_b I_bias_pos I_bias_neg VSS
*.PININFO V_LO:I V_LO_b:I V_RF:I V_RF_b:I V_out_p:O V_out_n:O I_bias_neg:B I_bias_pos:B VSS:B
M_LO_1_M1 V_out_p V_LO RF_M1_drain VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_LO_1_M2 V_out_n V_LO_b RF_M1_drain VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_LO_2_M1 V_out_p V_LO_b RF_M2_drain VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_LO_2_M2 V_out_n V_LO RF_M2_drain VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_RF_M1 RF_M1_drain V_RF I_bias_pos VSS nfet_03v3 L=0.28u W=10u nf=5 m=1
M_RF_M2 RF_M2_drain V_RF_b I_bias_neg VSS nfet_03v3 L=0.28u W=10u nf=5 m=1
M_RF_dummies VSS VSS VSS VSS nfet_03v3 L=0.28u W=2u nf=1 m=4
.ends
.end
