magic
tech gf180mcuD
magscale 1 10
timestamp 1757884110
<< pwell >>
rect -1176 -4524 1176 4524
<< mvpsubdiff >>
rect -1152 4487 1152 4500
rect -1152 4441 -1036 4487
rect 1036 4441 1152 4487
rect -1152 4428 1152 4441
rect -1152 4384 -1080 4428
rect -1152 2312 -1139 4384
rect -1093 2312 -1080 4384
rect 1080 4384 1152 4428
rect -1152 2268 -1080 2312
rect 1080 2312 1093 4384
rect 1139 2312 1152 4384
rect 1080 2268 1152 2312
rect -1152 2255 1152 2268
rect -1152 2209 -1036 2255
rect 1036 2209 1152 2255
rect -1152 2196 1152 2209
rect -1152 2152 -1080 2196
rect -1152 80 -1139 2152
rect -1093 80 -1080 2152
rect 1080 2152 1152 2196
rect -1152 36 -1080 80
rect 1080 80 1093 2152
rect 1139 80 1152 2152
rect 1080 36 1152 80
rect -1152 23 1152 36
rect -1152 -23 -1036 23
rect 1036 -23 1152 23
rect -1152 -36 1152 -23
rect -1152 -80 -1080 -36
rect -1152 -2152 -1139 -80
rect -1093 -2152 -1080 -80
rect 1080 -80 1152 -36
rect -1152 -2196 -1080 -2152
rect 1080 -2152 1093 -80
rect 1139 -2152 1152 -80
rect 1080 -2196 1152 -2152
rect -1152 -2209 1152 -2196
rect -1152 -2255 -1036 -2209
rect 1036 -2255 1152 -2209
rect -1152 -2268 1152 -2255
rect -1152 -2312 -1080 -2268
rect -1152 -4384 -1139 -2312
rect -1093 -4384 -1080 -2312
rect 1080 -2312 1152 -2268
rect -1152 -4428 -1080 -4384
rect 1080 -4384 1093 -2312
rect 1139 -4384 1152 -2312
rect 1080 -4428 1152 -4384
rect -1152 -4441 1152 -4428
rect -1152 -4487 -1036 -4441
rect 1036 -4487 1152 -4441
rect -1152 -4500 1152 -4487
<< mvpsubdiffcont >>
rect -1036 4441 1036 4487
rect -1139 2312 -1093 4384
rect 1093 2312 1139 4384
rect -1036 2209 1036 2255
rect -1139 80 -1093 2152
rect 1093 80 1139 2152
rect -1036 -23 1036 23
rect -1139 -2152 -1093 -80
rect 1093 -2152 1139 -80
rect -1036 -2255 1036 -2209
rect -1139 -4384 -1093 -2312
rect 1093 -4384 1139 -2312
rect -1036 -4487 1036 -4441
<< mvndiode >>
rect -1000 4335 1000 4348
rect -1000 2361 -987 4335
rect 987 2361 1000 4335
rect -1000 2348 1000 2361
rect -1000 2103 1000 2116
rect -1000 129 -987 2103
rect 987 129 1000 2103
rect -1000 116 1000 129
rect -1000 -129 1000 -116
rect -1000 -2103 -987 -129
rect 987 -2103 1000 -129
rect -1000 -2116 1000 -2103
rect -1000 -2361 1000 -2348
rect -1000 -4335 -987 -2361
rect 987 -4335 1000 -2361
rect -1000 -4348 1000 -4335
<< mvndiodec >>
rect -987 2361 987 4335
rect -987 129 987 2103
rect -987 -2103 987 -129
rect -987 -4335 987 -2361
<< metal1 >>
rect -1139 4441 -1036 4487
rect 1036 4441 1139 4487
rect -1139 4384 -1093 4441
rect 1093 4384 1139 4441
rect -998 2361 -987 4335
rect 987 2361 998 4335
rect -1139 2255 -1093 2312
rect 1093 2255 1139 2312
rect -1139 2209 -1036 2255
rect 1036 2209 1139 2255
rect -1139 2152 -1093 2209
rect 1093 2152 1139 2209
rect -998 129 -987 2103
rect 987 129 998 2103
rect -1139 23 -1093 80
rect 1093 23 1139 80
rect -1139 -23 -1036 23
rect 1036 -23 1139 23
rect -1139 -80 -1093 -23
rect 1093 -80 1139 -23
rect -998 -2103 -987 -129
rect 987 -2103 998 -129
rect -1139 -2209 -1093 -2152
rect 1093 -2209 1139 -2152
rect -1139 -2255 -1036 -2209
rect 1036 -2255 1139 -2209
rect -1139 -2312 -1093 -2255
rect 1093 -2312 1139 -2255
rect -998 -4335 -987 -2361
rect 987 -4335 998 -2361
rect -1139 -4441 -1093 -4384
rect 1093 -4441 1139 -4384
rect -1139 -4487 -1036 -4441
rect 1036 -4487 1139 -4441
<< properties >>
string diode_nd2ps_06v0_9F7MZ3 parameters
string FIXED_BBOX -1116 2232 1116 4464
string gencell diode_nd2ps_06v0
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 1 ny 4 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 doverlap 1 full_metal 1 compatible {diode_nd2ps_03v3 diode_nd2ps_06v0}
<< end >>
