magic
tech gf180mcuD
magscale 1 10
timestamp 1757961865
<< metal1 >>
rect 2599 10790 3478 10792
rect 2599 10787 7150 10790
rect -7273 10780 7150 10787
rect -7273 10362 7530 10780
rect -7273 10036 -6315 10362
rect 2390 10036 7530 10362
rect -7273 9982 7530 10036
rect 3350 9980 7530 9982
rect 2447 9698 2531 9700
rect -6424 9608 -6409 9698
rect 2508 9608 2531 9698
rect 2447 9602 2531 9608
rect -5943 7732 -5933 8316
rect -4592 7732 -4582 8316
rect -3726 7713 -3716 8297
rect -2375 7713 -2365 8297
rect -1501 7709 -1491 8293
rect -150 7709 -140 8293
rect 680 7723 690 8307
rect 2031 7723 2041 8307
rect 4170 6870 7530 9980
rect -6320 -810 2950 -800
rect -7200 -1620 2950 -810
rect -7200 -1650 -6360 -1620
rect 2500 -1650 2950 -1620
rect 4170 -1350 4630 6870
rect 4680 6760 4810 6770
rect 4680 -1230 4690 6760
rect 4800 -1230 4810 6760
rect 4680 -1240 4810 -1230
rect 6880 6760 7010 6770
rect 6880 -1230 6890 6760
rect 7000 -1230 7010 6760
rect 6880 -1240 7010 -1230
rect 7070 -1350 7530 6870
rect -7200 -3810 -6358 -1650
rect -5942 -2413 -5932 -1829
rect -4591 -2413 -4581 -1829
rect -3725 -2413 -3715 -1829
rect -2374 -2413 -2364 -1829
rect -1500 -2410 -1490 -1826
rect -149 -2410 -139 -1826
rect 680 -2410 690 -1826
rect 2031 -2410 2041 -1826
rect 2500 -1880 2952 -1650
rect 2502 -3810 2952 -1880
rect 4170 -2080 7530 -1350
rect -7200 -4830 2952 -3810
<< via1 >>
rect -6315 10036 2390 10362
rect -6409 9608 2508 9698
rect -5933 7732 -4592 8316
rect -3716 7713 -2375 8297
rect -1491 7709 -150 8293
rect 690 7723 2031 8307
rect 4690 -1230 4800 6760
rect 6890 -1230 7000 6760
rect -5932 -2413 -4591 -1829
rect -3715 -2413 -2374 -1829
rect -1490 -2410 -149 -1826
rect 690 -2410 2031 -1826
<< metal2 >>
rect -6433 10362 2539 10493
rect -6433 10036 -6315 10362
rect 2390 10036 2539 10362
rect -6433 9930 2539 10036
rect -6431 9698 2538 9930
rect -6431 9608 -6409 9698
rect 2508 9608 2538 9698
rect -6431 9595 2538 9608
rect -5950 8316 -4570 8330
rect -5950 7732 -5933 8316
rect -4592 7732 -4570 8316
rect -5950 6760 -4570 7732
rect -3730 8297 -2350 8330
rect -3730 7713 -3716 8297
rect -2375 7713 -2350 8297
rect -3730 6760 -2350 7713
rect -1510 8293 -130 8330
rect -1510 7709 -1491 8293
rect -150 7709 -130 8293
rect -1510 6760 -130 7709
rect 670 8307 2050 8320
rect 670 7723 690 8307
rect 2031 7723 2050 8307
rect 670 6770 2050 7723
rect 670 6760 4810 6770
rect -7220 -1230 4690 6760
rect 4800 -1230 4810 6760
rect -7220 -1240 4810 -1230
rect 6880 6760 7930 6770
rect 6880 -1230 6890 6760
rect 7000 -1230 7930 6760
rect 6880 -1240 7930 -1230
rect -5950 -1829 -4570 -1240
rect -5950 -2413 -5932 -1829
rect -4591 -2413 -4570 -1829
rect -5950 -2420 -4570 -2413
rect -3730 -1829 -2350 -1240
rect -3730 -2413 -3715 -1829
rect -2374 -2413 -2350 -1829
rect -3730 -2420 -2350 -2413
rect -1510 -1826 -130 -1240
rect -1510 -2410 -1490 -1826
rect -149 -2410 -130 -1826
rect -1510 -2420 -130 -2410
rect 670 -1826 2050 -1240
rect 670 -2410 690 -1826
rect 2031 -2410 2050 -1826
rect 670 -2430 2050 -2410
use diode_nd2ps_06v0_MV3SZ3  diode_nd2ps_06v0_MV3SZ3_0
timestamp 1757961865
transform 1 0 -1916 0 1 -2714
box -4524 -1176 4524 1176
use diode_pd2nw_06v0_5DG9HC  diode_pd2nw_06v0_5DG9HC_0
timestamp 1757961865
transform 1 0 -1944 0 1 8542
box -4676 -1352 4676 1352
use ppolyf_u_9H3LNU  ppolyf_u_9H3LNU_0
timestamp 1757961865
transform 0 1 5848 -1 0 2766
box -4216 -1318 4216 1318
<< labels >>
rlabel metal1 -7168 10450 -7168 10450 1 VDD
port 2 n
rlabel metal1 -6708 -4450 -6708 -4450 1 VSS
port 3 n
rlabel metal2 7740 3020 7740 3020 1 ASIG5V
port 0 n
rlabel metal2 -6710 3260 -6710 3280 1 to_gate
port 1 n
<< end >>
