magic
tech gf180mcuD
magscale 1 10
timestamp 1757884110
<< nwell >>
rect -616 -718 616 718
<< nsubdiff >>
rect -592 622 592 694
rect -592 578 -520 622
rect -592 -578 -579 578
rect -533 -578 -520 578
rect 520 578 592 622
rect -592 -622 -520 -578
rect 520 -578 533 578
rect 579 -578 592 578
rect 520 -622 592 -578
rect -592 -694 592 -622
<< nsubdiffcont >>
rect -579 -578 -533 578
rect 533 -578 579 578
<< polysilicon >>
rect -400 489 400 502
rect -400 443 -387 489
rect 387 443 400 489
rect -400 400 400 443
rect -400 -443 400 -400
rect -400 -489 -387 -443
rect 387 -489 400 -443
rect -400 -502 400 -489
<< polycontact >>
rect -387 443 387 489
rect -387 -489 387 -443
<< ppolyres >>
rect -400 -400 400 400
<< metal1 >>
rect -579 635 579 681
rect -579 578 -533 635
rect 533 578 579 635
rect -398 443 -387 489
rect 387 443 398 489
rect -398 -489 -387 -443
rect 387 -489 398 -443
rect -579 -635 -533 -578
rect 533 -635 579 -578
rect -579 -681 579 -635
<< properties >>
string FIXED_BBOX -556 -658 556 658
string gencell ppolyf_u
string library gf180mcu
string parameters w 4.0 l 4.0 m 1 nx 1 wmin 0.80 lmin 1.00 class resistor rho 315 val 320.61 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 1 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
string ppolyf_u_QK93DU parameters
<< end >>
