magic
tech gf180mcuD
magscale 1 10
timestamp 1757884110
<< nwell >>
rect -4803 -1176 4803 1176
<< pwell >>
rect -4979 1176 4979 1352
rect -4979 -1176 -4803 1176
rect 4803 -1176 4979 1176
rect -4979 -1352 4979 -1176
<< mvpsubdiff >>
rect -4947 1248 4947 1320
rect -4947 1204 -4875 1248
rect -4947 -1204 -4934 1204
rect -4888 -1204 -4875 1204
rect 4875 1204 4947 1248
rect -4947 -1248 -4875 -1204
rect 4875 -1204 4888 1204
rect 4934 -1204 4947 1204
rect 4875 -1248 4947 -1204
rect -4947 -1320 4947 -1248
<< mvnsubdiff >>
rect -4771 1131 -2483 1144
rect -4771 1085 -4655 1131
rect -2599 1085 -2483 1131
rect -4771 1072 -2483 1085
rect -4771 1028 -4699 1072
rect -4771 -1028 -4758 1028
rect -4712 -1028 -4699 1028
rect -2555 1028 -2483 1072
rect -4771 -1072 -4699 -1028
rect -2555 -1028 -2542 1028
rect -2496 -1028 -2483 1028
rect -2555 -1072 -2483 -1028
rect -4771 -1085 -2483 -1072
rect -4771 -1131 -4655 -1085
rect -2599 -1131 -2483 -1085
rect -4771 -1144 -2483 -1131
rect -2353 1131 -65 1144
rect -2353 1085 -2237 1131
rect -181 1085 -65 1131
rect -2353 1072 -65 1085
rect -2353 1028 -2281 1072
rect -2353 -1028 -2340 1028
rect -2294 -1028 -2281 1028
rect -137 1028 -65 1072
rect -2353 -1072 -2281 -1028
rect -137 -1028 -124 1028
rect -78 -1028 -65 1028
rect -137 -1072 -65 -1028
rect -2353 -1085 -65 -1072
rect -2353 -1131 -2237 -1085
rect -181 -1131 -65 -1085
rect -2353 -1144 -65 -1131
rect 65 1131 2353 1144
rect 65 1085 181 1131
rect 2237 1085 2353 1131
rect 65 1072 2353 1085
rect 65 1028 137 1072
rect 65 -1028 78 1028
rect 124 -1028 137 1028
rect 2281 1028 2353 1072
rect 65 -1072 137 -1028
rect 2281 -1028 2294 1028
rect 2340 -1028 2353 1028
rect 2281 -1072 2353 -1028
rect 65 -1085 2353 -1072
rect 65 -1131 181 -1085
rect 2237 -1131 2353 -1085
rect 65 -1144 2353 -1131
rect 2483 1131 4771 1144
rect 2483 1085 2599 1131
rect 4655 1085 4771 1131
rect 2483 1072 4771 1085
rect 2483 1028 2555 1072
rect 2483 -1028 2496 1028
rect 2542 -1028 2555 1028
rect 4699 1028 4771 1072
rect 2483 -1072 2555 -1028
rect 4699 -1028 4712 1028
rect 4758 -1028 4771 1028
rect 4699 -1072 4771 -1028
rect 2483 -1085 4771 -1072
rect 2483 -1131 2599 -1085
rect 4655 -1131 4771 -1085
rect 2483 -1144 4771 -1131
<< mvpsubdiffcont >>
rect -4934 -1204 -4888 1204
rect 4888 -1204 4934 1204
<< mvnsubdiffcont >>
rect -4655 1085 -2599 1131
rect -4758 -1028 -4712 1028
rect -2542 -1028 -2496 1028
rect -4655 -1131 -2599 -1085
rect -2237 1085 -181 1131
rect -2340 -1028 -2294 1028
rect -124 -1028 -78 1028
rect -2237 -1131 -181 -1085
rect 181 1085 2237 1131
rect 78 -1028 124 1028
rect 2294 -1028 2340 1028
rect 181 -1131 2237 -1085
rect 2599 1085 4655 1131
rect 2496 -1028 2542 1028
rect 4712 -1028 4758 1028
rect 2599 -1131 4655 -1085
<< mvpdiode >>
rect -4627 987 -2627 1000
rect -4627 -987 -4614 987
rect -2640 -987 -2627 987
rect -4627 -1000 -2627 -987
rect -2209 987 -209 1000
rect -2209 -987 -2196 987
rect -222 -987 -209 987
rect -2209 -1000 -209 -987
rect 209 987 2209 1000
rect 209 -987 222 987
rect 2196 -987 2209 987
rect 209 -1000 2209 -987
rect 2627 987 4627 1000
rect 2627 -987 2640 987
rect 4614 -987 4627 987
rect 2627 -1000 4627 -987
<< mvpdiodec >>
rect -4614 -987 -2640 987
rect -2196 -987 -222 987
rect 222 -987 2196 987
rect 2640 -987 4614 987
<< metal1 >>
rect -4934 1261 4934 1307
rect -4934 1204 -4888 1261
rect 4888 1204 4934 1261
rect -4758 1085 -4655 1131
rect -2599 1085 -2496 1131
rect -4758 1028 -4712 1085
rect -2542 1028 -2496 1085
rect -4625 -987 -4614 987
rect -2640 -987 -2629 987
rect -4758 -1085 -4712 -1028
rect -2542 -1085 -2496 -1028
rect -4758 -1131 -4655 -1085
rect -2599 -1131 -2496 -1085
rect -2340 1085 -2237 1131
rect -181 1085 -78 1131
rect -2340 1028 -2294 1085
rect -124 1028 -78 1085
rect -2207 -987 -2196 987
rect -222 -987 -211 987
rect -2340 -1085 -2294 -1028
rect -124 -1085 -78 -1028
rect -2340 -1131 -2237 -1085
rect -181 -1131 -78 -1085
rect 78 1085 181 1131
rect 2237 1085 2340 1131
rect 78 1028 124 1085
rect 2294 1028 2340 1085
rect 211 -987 222 987
rect 2196 -987 2207 987
rect 78 -1085 124 -1028
rect 2294 -1085 2340 -1028
rect 78 -1131 181 -1085
rect 2237 -1131 2340 -1085
rect 2496 1085 2599 1131
rect 4655 1085 4758 1131
rect 2496 1028 2542 1085
rect 4712 1028 4758 1085
rect 2629 -987 2640 987
rect 4614 -987 4625 987
rect 2496 -1085 2542 -1028
rect 4712 -1085 4758 -1028
rect 2496 -1131 2599 -1085
rect 4655 -1131 4758 -1085
rect -4934 -1261 -4888 -1204
rect 4888 -1261 4934 -1204
rect -4934 -1307 4934 -1261
<< properties >>
string diode_pd2nw_06v0_5DGPGC parameters
string FIXED_BBOX 2519 -1108 4735 1108
string gencell diode_pd2nw_06v0
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 4 ny 1 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 0 gbc 0 doverlap 0 full_metal 1 compatible {diode_pd2nw_03v3 diode_pd2nw_06v0}
<< end >>
