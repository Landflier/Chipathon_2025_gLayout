magic
tech gf180mcuD
magscale 1 10
timestamp 1757884110
<< pwell >>
rect -4524 -1176 4524 1176
<< mvpsubdiff >>
rect -4500 1139 4500 1152
rect -4500 1093 -4384 1139
rect -2312 1093 -2152 1139
rect -80 1093 80 1139
rect 2152 1093 2312 1139
rect 4384 1093 4500 1139
rect -4500 1080 4500 1093
rect -4500 1036 -4428 1080
rect -4500 -1036 -4487 1036
rect -4441 -1036 -4428 1036
rect -2268 1036 -2196 1080
rect -4500 -1080 -4428 -1036
rect -2268 -1036 -2255 1036
rect -2209 -1036 -2196 1036
rect -36 1036 36 1080
rect -2268 -1080 -2196 -1036
rect -36 -1036 -23 1036
rect 23 -1036 36 1036
rect 2196 1036 2268 1080
rect -36 -1080 36 -1036
rect 2196 -1036 2209 1036
rect 2255 -1036 2268 1036
rect 4428 1036 4500 1080
rect 2196 -1080 2268 -1036
rect 4428 -1036 4441 1036
rect 4487 -1036 4500 1036
rect 4428 -1080 4500 -1036
rect -4500 -1093 4500 -1080
rect -4500 -1139 -4384 -1093
rect -2312 -1139 -2152 -1093
rect -80 -1139 80 -1093
rect 2152 -1139 2312 -1093
rect 4384 -1139 4500 -1093
rect -4500 -1152 4500 -1139
<< mvpsubdiffcont >>
rect -4384 1093 -2312 1139
rect -2152 1093 -80 1139
rect 80 1093 2152 1139
rect 2312 1093 4384 1139
rect -4487 -1036 -4441 1036
rect -2255 -1036 -2209 1036
rect -23 -1036 23 1036
rect 2209 -1036 2255 1036
rect 4441 -1036 4487 1036
rect -4384 -1139 -2312 -1093
rect -2152 -1139 -80 -1093
rect 80 -1139 2152 -1093
rect 2312 -1139 4384 -1093
<< mvndiode >>
rect -4348 987 -2348 1000
rect -4348 -987 -4335 987
rect -2361 -987 -2348 987
rect -4348 -1000 -2348 -987
rect -2116 987 -116 1000
rect -2116 -987 -2103 987
rect -129 -987 -116 987
rect -2116 -1000 -116 -987
rect 116 987 2116 1000
rect 116 -987 129 987
rect 2103 -987 2116 987
rect 116 -1000 2116 -987
rect 2348 987 4348 1000
rect 2348 -987 2361 987
rect 4335 -987 4348 987
rect 2348 -1000 4348 -987
<< mvndiodec >>
rect -4335 -987 -2361 987
rect -2103 -987 -129 987
rect 129 -987 2103 987
rect 2361 -987 4335 987
<< metal1 >>
rect -4487 1093 -4384 1139
rect -2312 1093 -2152 1139
rect -80 1093 80 1139
rect 2152 1093 2312 1139
rect 4384 1093 4487 1139
rect -4487 1036 -4441 1093
rect -2255 1036 -2209 1093
rect -4346 -987 -4335 987
rect -2361 -987 -2350 987
rect -4487 -1093 -4441 -1036
rect -23 1036 23 1093
rect -2114 -987 -2103 987
rect -129 -987 -118 987
rect -2255 -1093 -2209 -1036
rect 2209 1036 2255 1093
rect 118 -987 129 987
rect 2103 -987 2114 987
rect -23 -1093 23 -1036
rect 4441 1036 4487 1093
rect 2350 -987 2361 987
rect 4335 -987 4346 987
rect 2209 -1093 2255 -1036
rect 4441 -1093 4487 -1036
rect -4487 -1139 -4384 -1093
rect -2312 -1139 -2152 -1093
rect -80 -1139 80 -1093
rect 2152 -1139 2312 -1093
rect 4384 -1139 4487 -1093
<< properties >>
string diode_nd2ps_06v0_MV3SZ3 parameters
string FIXED_BBOX 2232 -1116 4464 1116
string gencell diode_nd2ps_06v0
string library gf180mcu
string parameters w 10 l 10 area 100.0 peri 40.0 nx 4 ny 1 dummy 0 lmin 0.45 wmin 0.45 class diode elc 1 erc 1 etc 1 ebc 1 doverlap 1 full_metal 1 compatible {diode_nd2ps_03v3 diode_nd2ps_06v0}
<< end >>
