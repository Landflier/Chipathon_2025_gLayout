** sch_path: /home/vasil/Downloads/SSCS_PICO_2025/src/design_xsch/Gilbert_cell_no_hierarchy.sch
.subckt Gilbert_cell_no_hierarchy VDD V_out_p V_out_n V_LO V_LO_b V_RF V_RF_b I_bias_pos I_bias_neg VSS
*.PININFO V_LO:I V_LO_b:I V_RF:I V_RF_b:I V_out_p:O V_out_n:O I_bias_neg:B I_bias_pos:B VDD:B VSS:B
M_dp_lo_pos V_out_p V_LO rf_diff_pair_pos_input VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_dp_lo_neg V_out_n V_LO_b rf_diff_pair_pos_input VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_dp_lo_b_pos V_out_p V_LO_b rf_diff_pair_neg_input VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_dp_lo_b_neg V_out_n V_LO rf_diff_pair_neg_input VSS nfet_03v3 L=0.28u W=20u nf=5 m=1
M_rf_pos rf_diff_pair_pos_input V_RF I_bias_pos VSS nfet_03v3 L=0.28u W=10u nf=5 m=1
M_rf_neg rf_diff_pair_neg_input V_RF_b I_bias_neg VSS nfet_03v3 L=0.28u W=10u nf=5 m=1
XR_load_1 V_out_n VDD VSS pplus_u r_width=2e-6 r_length=10e-6 m=1
XR_load_2 V_out_p VDD VSS pplus_u r_width=2e-6 r_length=10e-6 m=1
XR_degen I_bias_neg I_bias_pos VSS pplus_u r_width=1e-6 r_length=7e-6 m=1
.ends
.end
