magic
tech gf180mcuD
magscale 1 5
timestamp 1755250493
<< checkpaint >>
rect -534 1090 1744 1120
rect -534 780 1992 1090
rect -1030 -2030 1992 780
rect -782 -2060 1992 -2030
rect -534 -2090 1992 -2060
rect -286 -2120 1992 -2090
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
use pfet_03v3_KAQ8RX  M1
timestamp 0
transform 1 0 605 0 1 -485
box -139 -605 139 605
use pfet_03v3_KAQ8RX  M2
timestamp 0
transform 1 0 853 0 1 -515
box -139 -605 139 605
use nfet_03v3_WYMPLR  M3
timestamp 0
transform 1 0 109 0 1 -625
box -139 -405 139 405
use nfet_03v3_WYMPLR  M4
timestamp 0
transform 1 0 357 0 1 -655
box -139 -405 139 405
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 Vout
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 Vin_plus
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 640 0 0 0 Vin_minus
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 640 0 0 0 I_bias
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 640 0 0 0 VSS
port 5 nsew
<< end >>
