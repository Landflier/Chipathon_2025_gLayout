magic
tech gf180mcuD
magscale 1 10
timestamp 1757925023
<< pwell >>
rect -6727 -6681 -6687 -4604
<< metal1 >>
rect -7650 -560 6280 110
rect -7650 -2680 -6880 -560
rect 2710 -1830 6280 -560
rect -6400 -2510 -6390 -2000
rect -5020 -2510 -5010 -2000
rect -4130 -2490 -4120 -1980
rect -2750 -2490 -2740 -1980
rect -1770 -2490 -1760 -1980
rect -390 -2490 -380 -1980
rect 590 -2500 600 -1990
rect 1970 -2500 1980 -1990
rect 2710 -2680 4610 -1830
rect -7650 -3320 4610 -2680
rect -7230 -4550 2470 -4160
rect -7230 -6451 -6735 -4550
rect -7230 -6690 -6733 -6451
rect -6637 -6627 -6627 -4653
rect -6390 -5350 -6380 -4840
rect -5010 -5350 -5000 -4840
rect -4653 -6627 -4643 -4653
rect -4120 -5300 -4110 -4790
rect -2740 -5300 -2730 -4790
rect -1760 -5310 -1750 -4800
rect -380 -5310 -370 -4800
rect 580 -5250 590 -4740
rect 1960 -5250 1970 -4740
rect 2134 -6690 2464 -4550
rect 3820 -5290 4610 -3320
rect 4670 -3280 4810 -3270
rect 4670 -4150 4700 -3280
rect 4800 -4150 4810 -3280
rect 4670 -4170 4810 -4150
rect 5650 -3280 5780 -3270
rect 5650 -4150 5660 -3280
rect 5760 -4150 5780 -3280
rect 5650 -4170 5780 -4150
rect 5860 -5290 6280 -1830
rect 3820 -5590 6280 -5290
rect -7230 -7349 2464 -6690
rect -7230 -7359 2450 -7349
rect -7230 -7360 -7150 -7359
rect -6622 -7360 2450 -7359
<< via1 >>
rect -6390 -2510 -5020 -2000
rect -4120 -2490 -2750 -1980
rect -1760 -2490 -390 -1980
rect 600 -2500 1970 -1990
rect -6380 -5350 -5010 -4840
rect -4110 -5300 -2740 -4790
rect -1750 -5310 -380 -4800
rect 590 -5250 1960 -4740
rect 4700 -4150 4800 -3280
rect 5660 -4150 5760 -3280
<< metal2 >>
rect -6430 -2000 -4994 -1888
rect -6430 -2510 -6390 -2000
rect -5020 -2510 -4994 -2000
rect -6430 -3250 -4994 -2510
rect -4150 -1980 -2714 -1828
rect -4150 -2490 -4120 -1980
rect -2750 -2490 -2714 -1980
rect -4150 -3250 -2714 -2490
rect -1790 -1980 -354 -1888
rect -1790 -2490 -1760 -1980
rect -390 -2490 -354 -1980
rect -1790 -3250 -354 -2490
rect 560 -1990 1996 -1928
rect 560 -2500 600 -1990
rect 1970 -2500 1996 -1990
rect 560 -3250 1996 -2500
rect -8160 -3280 4830 -3250
rect -8160 -4150 4700 -3280
rect 4800 -4150 4830 -3280
rect -8160 -4180 4830 -4150
rect 5650 -3280 6750 -3270
rect 5650 -4150 5660 -3280
rect 5760 -4150 6750 -3280
rect 5650 -4160 6750 -4150
rect -6430 -4643 -4994 -4180
rect -6627 -4653 -4653 -4643
rect -6430 -4840 -4994 -4653
rect -6430 -5350 -6380 -4840
rect -5010 -5350 -4994 -4840
rect -6430 -5520 -4994 -5350
rect -4150 -4790 -2714 -4180
rect -4150 -5300 -4110 -4790
rect -2740 -5300 -2714 -4790
rect -4150 -5460 -2714 -5300
rect -1790 -4800 -354 -4180
rect -1790 -5310 -1750 -4800
rect -380 -5310 -354 -4800
rect -1790 -5520 -354 -5310
rect 560 -4740 1996 -4180
rect 560 -5250 590 -4740
rect 1960 -5250 1996 -4740
rect 560 -5560 1996 -5250
rect -6627 -6637 -4653 -6627
<< rmetal2 >>
rect -6627 -5520 -6430 -4653
rect -4994 -5520 -4653 -4653
rect -6627 -6627 -4653 -5520
use diode_nd2ps_06v0_MV3SZ3  diode_nd2ps_06v0_MV3SZ3_0
timestamp 1757884110
transform 1 0 -2292 0 1 -5640
box -4524 -1176 4524 1176
use diode_pd2nw_06v0_5DGPGC  diode_pd2nw_06v0_5DGPGC_0
timestamp 1757884110
transform 1 0 -2181 0 1 -1608
box -4979 -1352 4979 1352
use ppolyf_u_4VJXJK  ppolyf_u_4VJXJK_0
timestamp 1757884110
transform 0 1 5228 -1 0 -3564
box -1816 -718 1816 718
<< labels >>
rlabel metal1 -7210 -5830 -7210 -5830 3 VSS
port 3 e
rlabel metal1 -7540 -1380 -7540 -1380 3 VDD
port 4 e
rlabel metal2 -7990 -3900 -7990 -3900 1 to_gate
port 5 n
rlabel metal2 6650 -3720 6650 -3720 1 ASIG5V
port 6 n
<< end >>
