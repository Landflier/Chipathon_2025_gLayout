* NGSPICE file created from nmos_Cmirror_with_decap_layout.ext - technology: gf180mcuD

.subckt Unnamed_278d0711 m4_n620_n620# m4_n500_n500# VSUBS
X0 m4_n500_n500# m4_n620_n620# cap_mim_2f0_m4m5_noshield c_width=5u c_length=5u
.ends

.subckt cmirror_interdigitized a_n2116_n809# a_n1852_n495# a_n1906_n75#
X0 a_n2116_n809# a_1322_n123# a_n1906_n75# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X1 a_n1906_n75# a_1622_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.855p pd=3.78u as=0.4575p ps=1.97u w=0.75u l=0.28u
X2 a_n1852_n495# a_n178_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X3 a_n2116_n809# a_n478_n123# a_n1906_n75# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X4 a_n1906_n75# a_n778_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X5 a_n2116_n809# a_n1078_n123# a_n1906_n75# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X6 a_n2116_n809# a_122_n123# a_n1852_n495# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X7 a_n1906_n75# a_n1378_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X8 a_n2116_n809# a_n1678_n123# a_n1906_n75# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.855p ps=3.78u w=0.75u l=0.28u
X9 a_n1906_n75# a_422_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X10 a_n2116_n809# a_722_n123# a_n1906_n75# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
X11 a_n1906_n75# a_1022_n123# a_n2116_n809# a_n2116_n809# nfet_03v3 ad=0.4575p pd=1.97u as=0.4575p ps=1.97u w=0.75u l=0.28u
.ends

.subckt nmos_Cmirror_with_decap_layout I_BIAS I_OUT VSS
XUnnamed_278d0711_0 I_BIAS VSS VSS Unnamed_278d0711
Xcmirror_interdigitized_0 VSS I_BIAS I_OUT cmirror_interdigitized
.ends

