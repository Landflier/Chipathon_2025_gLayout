magic
tech gf180mcuD
magscale 1 10
timestamp 1755084777
<< error_s >>
rect 1124 3203 1135 3249
rect 1181 3203 1192 3214
rect 1284 3203 1295 3249
rect 1341 3203 1352 3214
rect 1444 3203 1455 3249
rect 1501 3203 1512 3214
rect 1604 3203 1615 3249
rect 1661 3203 1672 3214
rect 1764 3203 1775 3249
rect 2684 3223 2695 3269
rect 2741 3223 2752 3234
rect 2844 3223 2855 3269
rect 2901 3223 2912 3234
rect 3004 3223 3015 3269
rect 3061 3223 3072 3234
rect 3164 3223 3175 3269
rect 3221 3223 3232 3234
rect 3324 3223 3335 3269
rect 3381 3223 3392 3234
rect 1821 3203 1832 3214
rect 4284 3203 4295 3249
rect 4341 3203 4352 3214
rect 4444 3203 4455 3249
rect 4501 3203 4512 3214
rect 4604 3203 4615 3249
rect 4661 3203 4672 3214
rect 4764 3203 4775 3249
rect 4821 3203 4832 3214
rect 4924 3203 4935 3249
rect 5794 3223 5805 3269
rect 5851 3223 5862 3234
rect 5954 3223 5965 3269
rect 6011 3223 6022 3234
rect 6114 3223 6125 3269
rect 6171 3223 6182 3234
rect 6274 3223 6285 3269
rect 6331 3223 6342 3234
rect 6434 3223 6445 3269
rect 6491 3223 6502 3234
rect 4981 3203 4992 3214
rect 2638 -808 2661 -797
rect 2775 -808 2821 -797
rect 2935 -808 2981 -797
rect 3095 -808 3141 -797
rect 3255 -808 3301 -797
rect 3415 -808 3438 -797
rect 5748 -808 5771 -797
rect 5885 -808 5931 -797
rect 6045 -808 6091 -797
rect 6205 -808 6251 -797
rect 6365 -808 6411 -797
rect 6525 -808 6548 -797
rect 1078 -828 1101 -817
rect 1215 -828 1261 -817
rect 1375 -828 1421 -817
rect 1535 -828 1581 -817
rect 1695 -828 1741 -817
rect 1855 -828 1878 -817
rect 4238 -828 4261 -817
rect 4375 -828 4421 -817
rect 4535 -828 4581 -817
rect 4695 -828 4741 -817
rect 4855 -828 4901 -817
rect 5015 -828 5038 -817
rect 1124 -909 1135 -863
rect 1284 -909 1295 -863
rect 1444 -909 1455 -863
rect 1604 -909 1615 -863
rect 1764 -909 1775 -863
rect 2684 -889 2695 -843
rect 2844 -889 2855 -843
rect 3004 -889 3015 -843
rect 3164 -889 3175 -843
rect 3324 -889 3335 -843
rect 4284 -909 4295 -863
rect 4444 -909 4455 -863
rect 4604 -909 4615 -863
rect 4764 -909 4775 -863
rect 4924 -909 4935 -863
rect 5794 -889 5805 -843
rect 5954 -889 5965 -843
rect 6114 -889 6125 -843
rect 6274 -889 6285 -843
rect 6434 -889 6445 -843
rect 1094 -1767 1105 -1721
rect 1151 -1767 1162 -1756
rect 1254 -1767 1265 -1721
rect 1311 -1767 1322 -1756
rect 1414 -1767 1425 -1721
rect 1471 -1767 1482 -1756
rect 1574 -1767 1585 -1721
rect 1631 -1767 1642 -1756
rect 1734 -1767 1745 -1721
rect 1791 -1767 1802 -1756
rect 2614 -1767 2625 -1721
rect 2671 -1767 2682 -1756
rect 2774 -1767 2785 -1721
rect 2831 -1767 2842 -1756
rect 2934 -1767 2945 -1721
rect 2991 -1767 3002 -1756
rect 3094 -1767 3105 -1721
rect 3151 -1767 3162 -1756
rect 3254 -1767 3265 -1721
rect 3311 -1767 3322 -1756
rect 1048 -3798 1071 -3787
rect 1185 -3798 1231 -3787
rect 1345 -3798 1391 -3787
rect 1505 -3798 1551 -3787
rect 1665 -3798 1711 -3787
rect 1825 -3798 1848 -3787
rect 2568 -3798 2591 -3787
rect 2705 -3798 2751 -3787
rect 2865 -3798 2911 -3787
rect 3025 -3798 3071 -3787
rect 3185 -3798 3231 -3787
rect 3345 -3798 3368 -3787
rect 1094 -3879 1105 -3833
rect 1254 -3879 1265 -3833
rect 1414 -3879 1425 -3833
rect 1574 -3879 1585 -3833
rect 1734 -3879 1745 -3833
rect 2614 -3879 2625 -3833
rect 2774 -3879 2785 -3833
rect 2934 -3879 2945 -3833
rect 3094 -3879 3105 -3833
rect 3254 -3879 3265 -3833
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use nfet_03v3_WQVELR  M_dp_lo_b_neg
timestamp 1755084777
transform 1 0 6148 0 1 1190
box -598 -2210 598 2210
use nfet_03v3_WQVELR  M_dp_lo_b_pos
timestamp 1755084777
transform 1 0 4638 0 1 1170
box -598 -2210 598 2210
use nfet_03v3_WQVELR  M_dp_lo_neg
timestamp 1755084777
transform 1 0 3038 0 1 1190
box -598 -2210 598 2210
use nfet_03v3_WQVELR  M_dp_lo_pos
timestamp 1755084777
transform 1 0 1478 0 1 1170
box -598 -2210 598 2210
use nfet_03v3_WQ9W9R  M_rf_neg
timestamp 1755084777
transform 1 0 2968 0 1 -2800
box -598 -1210 598 1210
use nfet_03v3_WQ9W9R  M_rf_pos
timestamp 1755084777
transform 1 0 1448 0 1 -2800
box -598 -1210 598 1210
use pplus_u_APHXDV  XR_degen
timestamp 1755084777
transform 1 0 6276 0 1 -2938
box -286 -1012 286 1012
use pplus_u_2PP5LV  XR_load_1
timestamp 1755084777
transform 1 0 4236 0 1 -2658
box -386 -1312 386 1312
use pplus_u_2PP5LV  XR_load_2
timestamp 1755084777
transform 1 0 5256 0 1 -2658
box -386 -1312 386 1312
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 1280 0 0 0 V_out_p
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 1280 0 0 0 V_out_n
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 1280 0 0 0 V_LO
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 1280 0 0 0 V_LO_b
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 1280 0 0 0 V_RF
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 1280 0 0 0 V_RF_b
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 1280 0 0 0 I_bias_pos
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 1280 0 0 0 I_bias_neg
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 1280 0 0 0 VSS
port 9 nsew
<< end >>
