magic
tech gf180mcuD
magscale 1 10
timestamp 1755084777
<< nwell >>
rect -286 -1012 286 1012
<< pdiff >>
rect -100 813 100 826
rect -100 767 -87 813
rect 87 767 100 813
rect -100 700 100 767
rect -100 -767 100 -700
rect -100 -813 -87 -767
rect 87 -813 100 -767
rect -100 -826 100 -813
<< pdiffc >>
rect -87 767 87 813
rect -87 -813 87 -767
<< nsubdiff >>
rect -262 916 262 988
rect -262 872 -190 916
rect -262 -872 -249 872
rect -203 -872 -190 872
rect 190 872 262 916
rect -262 -916 -190 -872
rect 190 -872 203 872
rect 249 -872 262 872
rect 190 -916 262 -872
rect -262 -988 262 -916
<< nsubdiffcont >>
rect -249 -872 -203 872
rect 203 -872 249 872
<< pdiffres >>
rect -100 -700 100 700
<< metal1 >>
rect -249 929 249 975
rect -249 872 -203 929
rect 203 872 249 929
rect -98 767 -87 813
rect 87 767 98 813
rect -98 -813 -87 -767
rect 87 -813 98 -767
rect -249 -929 -203 -872
rect 203 -929 249 -872
rect -249 -975 249 -929
<< properties >>
string FIXED_BBOX -226 -952 226 952
string gencell pplus_u
string library gf180mcu
string parameters w 1.0 l 7.0 m 1 nx 1 wmin 1.00 lmin 1.00 class resistor rho 128 val 914.285 dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.60 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
