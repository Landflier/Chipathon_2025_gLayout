magic
tech gf180mcuD
magscale 1 5
timestamp 1755250494
<< checkpaint >>
rect -286 1280 1992 1890
rect -1030 -1630 1992 1280
rect -782 -1660 1992 -1630
rect -534 -1690 1992 -1660
rect -286 -1720 1992 -1690
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
use nfet_03v3_WQ7QLR  M1
timestamp 0
transform 1 0 109 0 1 -175
box -139 -455 139 455
use nfet_03v3_VLS3DR  M2
timestamp 0
transform 1 0 357 0 1 -380
box -139 -280 139 280
use nfet_03v3_WQ7QLR  M3
timestamp 0
transform 1 0 605 0 1 -235
box -139 -455 139 455
use nfet_03v3_WG8W9R  M4
timestamp 0
transform 1 0 853 0 1 85
box -139 -805 139 805
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 I_BIAS
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 I_out_2
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 I_out_3
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 640 0 0 0 I_out_1
port 3 nsew
<< end >>
