magic
tech gf180mcuD
magscale 1 10
timestamp 1757869051
<< pwell >>
rect 550 430 2130 780
rect 550 410 1550 430
rect 550 180 1520 410
rect 1540 210 1720 390
rect 1570 180 1700 210
rect 1750 180 2130 430
rect 550 20 2130 180
rect 1570 -1120 1700 20
<< psubdiff >>
rect 550 410 2130 780
rect 550 180 1520 410
rect 1750 180 2130 410
rect 550 20 2130 180
<< ndiode >>
rect 1590 327 1680 340
rect 1590 263 1603 327
rect 1667 263 1680 327
rect 1590 250 1680 263
<< ndiodec >>
rect 1603 263 1667 327
<< metal1 >>
rect 550 410 2130 780
rect 550 180 1520 410
rect 1580 327 1690 350
rect 1580 263 1603 327
rect 1667 263 1690 327
rect 1580 240 1690 263
rect 1750 180 2130 410
rect 550 20 2130 180
rect 550 -430 750 -230
rect 4080 -420 4280 -220
rect 560 -950 2050 -660
rect 560 -1160 1520 -950
rect 1580 -1110 1690 -1000
rect 1750 -1160 2050 -950
rect 560 -1590 2050 -1160
<< metal2 >>
rect 1580 360 1690 370
rect 1580 220 1690 230
rect 750 -170 1760 -160
rect 750 -430 1560 -170
rect 1710 -430 1760 -170
rect 750 -440 1760 -430
rect 1580 -990 1690 -980
rect 1580 -1130 1690 -1120
<< via2 >>
rect 1580 230 1690 360
rect 1560 -430 1710 -170
rect 1580 -1120 1690 -990
<< metal3 >>
rect 1570 230 1580 360
rect 1690 230 1700 360
rect 1570 -170 1700 230
rect 1550 -430 1560 -170
rect 1710 -430 1720 -170
rect 1570 -990 1700 -430
rect 1570 -1120 1580 -990
rect 1690 -1120 1700 -990
use diode_nd2ps_03v3_A8G3GU  D1
timestamp 1757866917
transform 1 0 1635 0 1 -1055
box -205 -205 205 205
use diode_nd2ps_03v3_A8G3GU  D2
timestamp 1757866917
transform 1 0 1635 0 1 295
box -205 -205 205 205
use ppolyf_u_TZ73VR  XR1
timestamp 1757866917
transform 0 1 2898 -1 0 -324
box -316 -718 316 718
<< labels >>
flabel metal1 550 580 750 780 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 4080 -420 4280 -220 0 FreeSans 1280 0 0 0 ASIG5V
port 3 nsew
flabel metal1 550 -430 750 -230 0 FreeSans 1280 0 0 0 to_gate
port 1 nsew
flabel metal1 570 -1580 770 -1380 0 FreeSans 1280 0 0 0 VSS
port 2 nsew
<< end >>
