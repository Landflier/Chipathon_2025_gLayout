** sch_path: /home/vasil/Downloads/SSCS_PICO_2025/src/design_xsch/CMD_ESD_prot.sch
.subckt CMD_ESD_prot VDD to_gate VSS ASIG5V
*.PININFO VDD:B to_gate:B VSS:B ASIG5V:B
XR1 to_gate ASIG5V VDD ppolyf_u r_width=16e-6 r_length=4e-6 m=1
D1 to_gate VDD diode_pd2nw_06v0 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
D2 VSS to_gate diode_nd2ps_06v0 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
.ends
.end
