magic
tech gf180mcuD
magscale 1 5
timestamp 1755250493
<< checkpaint >>
rect -1030 2150 1248 2180
rect -1030 2120 1496 2150
rect -1030 2090 1744 2120
rect -1030 2060 1992 2090
rect -1030 2030 2240 2060
rect -1030 2000 2488 2030
rect -1030 -1030 2736 2000
rect -782 -1060 2736 -1030
rect -534 -1090 2736 -1060
rect -286 -1120 2736 -1090
rect -38 -1150 2736 -1120
rect 210 -1180 2736 -1150
rect 458 -1210 2736 -1180
<< metal1 >>
rect 0 0 100 100
use nfet_03v3_WG72DR  M_dummy_1
timestamp 0
transform 1 0 109 0 1 575
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_2
timestamp 0
transform 1 0 357 0 1 545
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_3
timestamp 0
transform 1 0 605 0 1 515
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_4
timestamp 0
transform 1 0 853 0 1 485
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_5
timestamp 0
transform 1 0 1101 0 1 455
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_6
timestamp 0
transform 1 0 1349 0 1 425
box -139 -605 139 605
use nfet_03v3_WG72DR  M_dummy_7
timestamp 0
transform 1 0 1597 0 1 395
box -139 -605 139 605
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 VSS
port 0 nsew
<< end >>
