magic
tech gf180mcuD
magscale 1 10
timestamp 1755084777
<< error_p >>
rect -354 1033 -343 1079
rect -297 1033 -286 1044
rect -194 1033 -183 1079
rect -137 1033 -126 1044
rect -34 1033 -23 1079
rect 23 1033 34 1044
rect 126 1033 137 1079
rect 183 1033 194 1044
rect 286 1033 297 1079
rect 343 1033 354 1044
rect -400 -998 -377 -987
rect -263 -998 -217 -987
rect -103 -998 -57 -987
rect 57 -998 103 -987
rect 217 -998 263 -987
rect 377 -998 400 -987
rect -354 -1079 -343 -1033
rect -194 -1079 -183 -1033
rect -34 -1079 -23 -1033
rect 126 -1079 137 -1033
rect 286 -1079 297 -1033
<< pwell >>
rect -598 -1210 598 1210
<< nmos >>
rect -348 -1000 -292 1000
rect -188 -1000 -132 1000
rect -28 -1000 28 1000
rect 132 -1000 188 1000
rect 292 -1000 348 1000
<< ndiff >>
rect -436 987 -348 1000
rect -436 -987 -423 987
rect -377 -987 -348 987
rect -436 -1000 -348 -987
rect -292 987 -188 1000
rect -292 -987 -263 987
rect -217 -987 -188 987
rect -292 -1000 -188 -987
rect -132 987 -28 1000
rect -132 -987 -103 987
rect -57 -987 -28 987
rect -132 -1000 -28 -987
rect 28 987 132 1000
rect 28 -987 57 987
rect 103 -987 132 987
rect 28 -1000 132 -987
rect 188 987 292 1000
rect 188 -987 217 987
rect 263 -987 292 987
rect 188 -1000 292 -987
rect 348 987 436 1000
rect 348 -987 377 987
rect 423 -987 436 987
rect 348 -1000 436 -987
<< ndiffc >>
rect -423 -987 -377 987
rect -263 -987 -217 987
rect -103 -987 -57 987
rect 57 -987 103 987
rect 217 -987 263 987
rect 377 -987 423 987
<< psubdiff >>
rect -574 1114 574 1186
rect -574 1070 -502 1114
rect -574 -1070 -561 1070
rect -515 -1070 -502 1070
rect 502 1070 574 1114
rect -574 -1114 -502 -1070
rect 502 -1070 515 1070
rect 561 -1070 574 1070
rect 502 -1114 574 -1070
rect -574 -1186 574 -1114
<< psubdiffcont >>
rect -561 -1070 -515 1070
rect 515 -1070 561 1070
<< polysilicon >>
rect -356 1079 -284 1092
rect -356 1033 -343 1079
rect -297 1033 -284 1079
rect -356 1020 -284 1033
rect -196 1079 -124 1092
rect -196 1033 -183 1079
rect -137 1033 -124 1079
rect -196 1020 -124 1033
rect -36 1079 36 1092
rect -36 1033 -23 1079
rect 23 1033 36 1079
rect -36 1020 36 1033
rect 124 1079 196 1092
rect 124 1033 137 1079
rect 183 1033 196 1079
rect 124 1020 196 1033
rect 284 1079 356 1092
rect 284 1033 297 1079
rect 343 1033 356 1079
rect 284 1020 356 1033
rect -348 1000 -292 1020
rect -188 1000 -132 1020
rect -28 1000 28 1020
rect 132 1000 188 1020
rect 292 1000 348 1020
rect -348 -1020 -292 -1000
rect -188 -1020 -132 -1000
rect -28 -1020 28 -1000
rect 132 -1020 188 -1000
rect 292 -1020 348 -1000
rect -356 -1033 -284 -1020
rect -356 -1079 -343 -1033
rect -297 -1079 -284 -1033
rect -356 -1092 -284 -1079
rect -196 -1033 -124 -1020
rect -196 -1079 -183 -1033
rect -137 -1079 -124 -1033
rect -196 -1092 -124 -1079
rect -36 -1033 36 -1020
rect -36 -1079 -23 -1033
rect 23 -1079 36 -1033
rect -36 -1092 36 -1079
rect 124 -1033 196 -1020
rect 124 -1079 137 -1033
rect 183 -1079 196 -1033
rect 124 -1092 196 -1079
rect 284 -1033 356 -1020
rect 284 -1079 297 -1033
rect 343 -1079 356 -1033
rect 284 -1092 356 -1079
<< polycontact >>
rect -343 1033 -297 1079
rect -183 1033 -137 1079
rect -23 1033 23 1079
rect 137 1033 183 1079
rect 297 1033 343 1079
rect -343 -1079 -297 -1033
rect -183 -1079 -137 -1033
rect -23 -1079 23 -1033
rect 137 -1079 183 -1033
rect 297 -1079 343 -1033
<< metal1 >>
rect -561 1127 561 1173
rect -561 1070 -515 1127
rect -354 1033 -343 1079
rect -297 1033 -286 1079
rect -194 1033 -183 1079
rect -137 1033 -126 1079
rect -34 1033 -23 1079
rect 23 1033 34 1079
rect 126 1033 137 1079
rect 183 1033 194 1079
rect 286 1033 297 1079
rect 343 1033 354 1079
rect 515 1070 561 1127
rect -423 987 -377 998
rect -423 -998 -377 -987
rect -263 987 -217 998
rect -263 -998 -217 -987
rect -103 987 -57 998
rect -103 -998 -57 -987
rect 57 987 103 998
rect 57 -998 103 -987
rect 217 987 263 998
rect 217 -998 263 -987
rect 377 987 423 998
rect 377 -998 423 -987
rect -561 -1127 -515 -1070
rect -354 -1079 -343 -1033
rect -297 -1079 -286 -1033
rect -194 -1079 -183 -1033
rect -137 -1079 -126 -1033
rect -34 -1079 -23 -1033
rect 23 -1079 34 -1033
rect 126 -1079 137 -1033
rect 183 -1079 194 -1033
rect 286 -1079 297 -1033
rect 343 -1079 354 -1033
rect 515 -1127 561 -1070
rect -561 -1173 561 -1127
<< properties >>
string FIXED_BBOX -538 -1150 538 1150
string gencell nfet_03v3
string library gf180mcu
string parameters w 10.0 l 0.28 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
